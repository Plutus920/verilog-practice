module jfkk(	input j,
		input k,		
		output q);
begin
